`ifndef UCODE_CTRL_VH_
`define UCODE_CTRL_VH_
`define INSTR_CTRL_SIZE 55
`define UCODE_ROM_SIZE 136

`define RESET_UCODE_INDEX 8'd128

`define INSTR_CTRL_SIGNALS_INDICES {6'd0, 6'd24, 6'd0, 6'd0, 6'd0, 6'd24, 6'd16, 6'd0, 6'd46, 6'd24, 6'd15, 6'd0, 6'd0, 6'd24, 6'd16, 6'd0, 6'd35, 6'd24, 6'd0, 6'd0, 6'd0, 6'd24, 6'd16, 6'd0, 6'd51, 6'd24, 6'd0, 6'd0, 6'd0, 6'd24, 6'd16, 6'd0, 6'd0, 6'd23, 6'd0, 6'd0, 6'd29, 6'd23, 6'd20, 6'd0, 6'd47, 6'd23, 6'd19, 6'd0, 6'd29, 6'd23, 6'd20, 6'd0, 6'd33, 6'd23, 6'd0, 6'd0, 6'd0, 6'd23, 6'd20, 6'd0, 6'd48, 6'd23, 6'd0, 6'd0, 6'd0, 6'd23, 6'd20, 6'd0, 6'd0, 6'd25, 6'd0, 6'd0, 6'd0, 6'd25, 6'd18, 6'd0, 6'd44, 6'd25, 6'd17, 6'd0, 6'd0, 6'd25, 6'd18, 6'd0, 6'd36, 6'd25, 6'd0, 6'd0, 6'd0, 6'd25, 6'd18, 6'd0, 6'd53, 6'd25, 6'd0, 6'd0, 6'd0, 6'd25, 6'd18, 6'd0, 6'd0, 6'd7, 6'd0, 6'd0, 6'd0, 6'd7, 6'd22, 6'd0, 6'd45, 6'd7, 6'd21, 6'd0, 6'd0, 6'd7, 6'd22, 6'd0, 6'd37, 6'd7, 6'd0, 6'd0, 6'd0, 6'd7, 6'd22, 6'd0, 6'd50, 6'd7, 6'd0, 6'd0, 6'd0, 6'd7, 6'd22, 6'd0, 6'd0, 6'd4, 6'd0, 6'd0, 6'd6, 6'd4, 6'd5, 6'd0, 6'd14, 6'd0, 6'd39, 6'd0, 6'd6, 6'd4, 6'd5, 6'd0, 6'd30, 6'd4, 6'd0, 6'd0, 6'd6, 6'd4, 6'd5, 6'd0, 6'd41, 6'd4, 6'd43, 6'd0, 6'd0, 6'd4, 6'd0, 6'd0, 6'd3, 6'd1, 6'd2, 6'd0, 6'd3, 6'd1, 6'd2, 6'd0, 6'd40, 6'd1, 6'd38, 6'd0, 6'd3, 6'd1, 6'd2, 6'd0, 6'd31, 6'd1, 6'd0, 6'd0, 6'd3, 6'd1, 6'd2, 6'd0, 6'd54, 6'd1, 6'd42, 6'd0, 6'd3, 6'd1, 6'd2, 6'd0, 6'd28, 6'd26, 6'd0, 6'd0, 6'd28, 6'd26, 6'd12, 6'd0, 6'd11, 6'd26, 6'd13, 6'd0, 6'd28, 6'd26, 6'd12, 6'd0, 6'd34, 6'd26, 6'd0, 6'd0, 6'd0, 6'd26, 6'd12, 6'd0, 6'd52, 6'd26, 6'd0, 6'd0, 6'd0, 6'd26, 6'd12, 6'd0, 6'd27, 6'd8, 6'd0, 6'd0, 6'd27, 6'd8, 6'd9, 6'd0, 6'd10, 6'd8, 6'd0, 6'd0, 6'd27, 6'd8, 6'd9, 6'd0, 6'd32, 6'd8, 6'd0, 6'd0, 6'd0, 6'd8, 6'd9, 6'd0, 6'd49, 6'd8, 6'd0, 6'd0, 6'd0, 6'd8, 6'd9, 6'd0}

`define INSTR_CTRL_SIGNALS_ROM {{ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_A, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_X, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_Y, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_X}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_Y}, {ALUOP_ADD, ALUDST_A, SRC1_A, SRC2_RMEM, 1'b0, ALUC_C, FLAG_ALU, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_A, SRC1_A, SRC2_RMEM, 1'b1, ALUC_C, FLAG_ALU, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b0, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_X, SRC1_X, SRC2_0, 1'b0, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_Y, SRC1_Y, SRC2_0, 1'b0, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b1, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_X, SRC1_X, SRC2_0, 1'b1, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_Y, SRC1_Y, SRC2_0, 1'b1, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_LEFT, ALUDST_A, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_LEFT, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_RIGHT, ALUDST_A, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_RIGHT, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_LEFT, ALUDST_A, SRC1_A, SRC2_0, 1'b0, ALUC_C, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_LEFT, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b0, ALUC_C, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_RIGHT, ALUDST_A, SRC1_A, SRC2_0, 1'b0, ALUC_C, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_SHIFT_RIGHT, ALUDST_WMEM, SRC1_RMEM, SRC2_0, 1'b0, ALUC_C, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_AND, ALUDST_A, SRC1_A, SRC2_RMEM, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_OR, ALUDST_A, SRC1_A, SRC2_RMEM, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_XOR, ALUDST_A, SRC1_A, SRC2_RMEM, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_NONE, SRC1_A, SRC2_RMEM, 1'b1, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_NONE, SRC1_X, SRC2_RMEM, 1'b1, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_NONE, SRC1_Y, SRC2_RMEM, 1'b1, ALUC_1, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_ALU, BRANCH_C, 1'b0, STORE_A}, {ALUOP_AND, ALUDST_NONE, SRC1_A, SRC2_RMEM, 1'b0, ALUC_0, FLAG_RMEM_BUFFER, FLAG_RMEM_BUFFER, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b1, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_Z, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_N, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_Z, 1'b1, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_N, 1'b1, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_V, 1'b1, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_V, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_X, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_A, SRC1_X, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_Y, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_A, SRC1_Y, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_X, SRC1_SP, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_SP, SRC1_X, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_ADD, ALUDST_A, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_ALU, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_ALU, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_STATUS}, {ALUOP_ADD, ALUDST_STATUS, SRC1_RMEM, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_1, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_1, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_1, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_0, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_0, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}, {ALUOP_HOLD, ALUDST_NONE, SRC1_A, SRC2_0, 1'b0, ALUC_0, FLAG_NONE, FLAG_0, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, FLAG_NONE, BRANCH_C, 1'b0, STORE_A}}

`define UCODE_CTRL_SIGNALS_INDICES {8'd1, 8'd92, 8'd0, 8'd0, 8'd0, 8'd45, 8'd48, 8'd0, 8'd16, 8'd31, 8'd29, 8'd0, 8'd0, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0, 8'd22, 8'd92, 8'd0, 8'd0, 8'd45, 8'd45, 8'd48, 8'd0, 8'd18, 8'd31, 8'd29, 8'd0, 8'd35, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0, 8'd7, 8'd92, 8'd0, 8'd0, 8'd0, 8'd45, 8'd48, 8'd0, 8'd16, 8'd31, 8'd29, 8'd0, 8'd33, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0, 8'd12, 8'd92, 8'd0, 8'd0, 8'd0, 8'd45, 8'd48, 8'd0, 8'd18, 8'd31, 8'd29, 8'd0, 8'd124, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0, 8'd0, 8'd104, 8'd0, 8'd0, 8'd51, 8'd51, 8'd51, 8'd0, 8'd27, 8'd0, 8'd27, 8'd0, 8'd43, 8'd43, 8'd43, 8'd0, 8'd89, 8'd120, 8'd0, 8'd0, 8'd64, 8'd64, 8'd66, 8'd0, 8'd27, 8'd86, 8'd27, 8'd0, 8'd0, 8'd83, 8'd0, 8'd0, 8'd31, 8'd92, 8'd31, 8'd0, 8'd45, 8'd45, 8'd45, 8'd0, 8'd27, 8'd31, 8'd27, 8'd0, 8'd35, 8'd35, 8'd35, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd52, 8'd52, 8'd56, 8'd0, 8'd27, 8'd73, 8'd27, 8'd0, 8'd68, 8'd68, 8'd73, 8'd0, 8'd31, 8'd92, 8'd0, 8'd0, 8'd45, 8'd45, 8'd48, 8'd0, 8'd27, 8'd31, 8'd27, 8'd0, 8'd35, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0, 8'd31, 8'd92, 8'd0, 8'd0, 8'd45, 8'd45, 8'd48, 8'd0, 8'd27, 8'd31, 8'd27, 8'd0, 8'd35, 8'd35, 8'd39, 8'd0, 8'd89, 8'd108, 8'd0, 8'd0, 8'd0, 8'd52, 8'd60, 8'd0, 8'd27, 8'd73, 8'd0, 8'd0, 8'd0, 8'd68, 8'd78, 8'd0}

`define UCODE_CTRL_SIGNALS_ROM {{ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_W, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_W, WMEMSRC_PCLO, SRC1_ALUOUT, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_W, WMEMSRC_STATUS_BRK, SRC1_ALUOUT, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_BRKLO, ADDRHI_FF, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_BRKHI, ADDRHI_FF, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_RMEM, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_PCLO, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_SP, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_SP, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_SP, ADDRHI_1, READ_EN_W, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_1, READ_EN_W, WMEMSRC_PCLO, SRC1_ALUOUT, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_RMEM_BUFFER, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b1, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b1, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_PCLO, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_BRANCH_BIT, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_BRANCH_BIT, 1'b0, BRANCH_DEPEND_BRANCH_BIT}, {ADDRLO_ALUOUT, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_PCHI, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_ALUOUT, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_NOT_C_OUT, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_NOT_C_OUT, 1'b0, BRANCH_DEPEND_NOT_C_OUT}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_ALUOUT, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_1, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_X, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_ALUOUT, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b1, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_RMEM, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_1, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_W, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_2, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_RMEM, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_0, READ_EN_R, WMEMSRC_PCHI, SRC1_Y, SRC2_RMEM, 1'b0, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_ALUCOUT, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_ALUOUT, READ_EN_W, WMEMSRC_INSTR_STORE, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_RMEM, SRC2_0, 1'b0, ALUC_1, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_1, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_RMEMBUFFER, ADDRHI_RMEM, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_ALUOUT, ADDRHI_HOLD, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_RMEM, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}, {ADDRLO_PCLO, ADDRHI_PCHI, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_SP, ADDRHI_1, READ_EN_R, WMEMSRC_PCHI, SRC1_SP, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_R, WMEMSRC_PCLO, SRC1_ALUOUT, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_R, WMEMSRC_STATUS_BC, SRC1_ALUOUT, SRC2_0, 1'b1, ALUC_0, ALUOP_ADD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_FC, ADDRHI_FF, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_ALUOUT, PCLOSRC_NONE, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_FD, ADDRHI_FF, READ_EN_R, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_RMEM, PCHISRC_NONE, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b1, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_0}, {ADDRLO_HOLD, ADDRHI_HOLD, READ_EN_NONE, WMEMSRC_PCHI, SRC1_A, SRC2_0, 1'b0, ALUC_0, ALUOP_HOLD, SPSRC_NONE, PCLOSRC_NONE, PCHISRC_RMEM, STATUS_SRC_NONE, BRANCH_DEPEND_0, INSTR_CTRL_0, 1'b0, BRANCH_DEPEND_0, 1'b0, BRANCH_DEPEND_1}}

`define DECODE_CTRL_SIGNALS_ROM {2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 2'd2, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd0, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd2, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd3, 2'd1, 2'd3, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd3, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd3, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0}

`endif