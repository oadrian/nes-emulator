
`define SAVE_STATE_BITS ($clog2(5080))

`define SAVE_STATE_LAST_ADDRESS 5080

`define SAVE_STATE_CPU_UCODE_INDEX 0
`define SAVE_STATE_CPU_INSTR_CTRL_INDEX 1
`define SAVE_STATE_CPU_STATE 2
`define SAVE_STATE_CPU_NMI_ACTIVE 3
`define SAVE_STATE_CPU_RESET_ACTIVE 4
`define SAVE_STATE_CPU_CURRENT_INTERRUPT 5
`define SAVE_STATE_CPU_A 6
`define SAVE_STATE_CPU_X 7
`define SAVE_STATE_CPU_Y 8
`define SAVE_STATE_CPU_SP 9
`define SAVE_STATE_CPU_N_FLAG 10
`define SAVE_STATE_CPU_V_FLAG 11
`define SAVE_STATE_CPU_D_FLAG 12
`define SAVE_STATE_CPU_I_FLAG 13
`define SAVE_STATE_CPU_Z_FLAG 14
`define SAVE_STATE_CPU_C_FLAG 15
`define SAVE_STATE_CPU_PC 16
`define SAVE_STATE_CPU_R_DATA_BUFFER 17
`define SAVE_STATE_CPU_ADDR 18
`define SAVE_STATE_CPU_ALU_OUT 19
`define SAVE_STATE_CPU_ALU_C_OUT 20
`define SAVE_STATE_CPU_ALU_V_OUT 21
`define SAVE_STATE_CPU_ALU_Z_OUT 22
`define SAVE_STATE_CPU_ALU_N_OUT 23
`define SAVE_STATE_CPU_MEM_CPU_RAM_LO 24
`define SAVE_STATE_CPU_MEM_CPU_RAM_HI 2071
`define SAVE_STATE_CPU_MEM_READ_DATA 2072
`define SAVE_STATE_CPU_MEM_PREV_REG_EN 2073
`define SAVE_STATE_CPU_MEM_PREV_BUT_RD 2074
`define SAVE_STATE_CPU_MEM_PREV_APU_RD 2075
`define SAVE_STATE_PPU_ROW 2076
`define SAVE_STATE_PPU_COL 2077
`define SAVE_STATE_PPU_HS_CURR_STATE 2078
`define SAVE_STATE_PPU_VS_CURR_STATE 2079
`define SAVE_STATE_PPU_PPU_BUF_IDX 2080
`define SAVE_STATE_PPU_PPU_BUFFER_LO 2081
`define SAVE_STATE_PPU_PPU_BUFFER_HI 2336
`define SAVE_STATE_PPU_VGA_BUFFER_LO 2337
`define SAVE_STATE_PPU_VGA_BUFFER_HI 2592
`define SAVE_STATE_PPU_TEMP_OAM_LO 2593
`define SAVE_STATE_PPU_TEMP_OAM_HI 2632
`define SAVE_STATE_PPU_TEMP_OAM_WR_IDX 2633
`define SAVE_STATE_PPU_TEMP_OAM_CNT 2634
`define SAVE_STATE_PPU_SEC_OAM_LO 2635
`define SAVE_STATE_PPU_SEC_OAM_HI 2674
`define SAVE_STATE_PPU_SEC_OAM_WR_IDX 2675
`define SAVE_STATE_PPU_SEC_OAM_CNT 2676
`define SAVE_STATE_REG_INTER_PPUCTRL_OUT 2677
`define SAVE_STATE_REG_INTER_PPUMASK_OUT 2678
`define SAVE_STATE_REG_INTER_OAMDMA_OUT 2679
`define SAVE_STATE_REG_INTER_OAMADDR_OUT 2680
`define SAVE_STATE_REG_INTER_WR_CURR_STATE 2681
`define SAVE_STATE_REG_INTER_REGDATA_OUT 2682
`define SAVE_STATE_REG_INTER_READ_BUF_CURR 2683
`define SAVE_STATE_REG_INTER_PPUSTATUS_OUT 2684
`define SAVE_STATE_REG_INTER_FORCE_VBLANK_CLR0 2685
`define SAVE_STATE_REG_INTER_FORCE_VBLANK_CLR1 2686
`define SAVE_STATE_REG_INTER_OAMDMA_CURR_STATE 2687
`define SAVE_STATE_REG_INTER_COUNTER 2688
`define SAVE_STATE_REG_INTER_FX 2689
`define SAVE_STATE_REG_INTER_TADDR 2690
`define SAVE_STATE_REG_INTER_VADDR 2691
`define SAVE_STATE_BG_PIXEL_NT 2692
`define SAVE_STATE_BG_PIXEL_AT 2693
`define SAVE_STATE_BG_PIXEL_BG_L 2694
`define SAVE_STATE_BG_PIXEL_BG_H 2695
`define SAVE_STATE_BG_PIXEL_BG_L_BOTH 2696
`define SAVE_STATE_BG_PIXEL_BG_H_BOTH 2697
`define SAVE_STATE_BG_PIXEL_AT_L_BOTH 2698
`define SAVE_STATE_BG_PIXEL_AT_H_BOTH 2699
`define SAVE_STATE_SP_EVAL_CURR_SPRITE 2700
`define SAVE_STATE_VGA_ROW_LO 2701
`define SAVE_STATE_VGA_ROW_HI 2710
`define SAVE_STATE_VGA_COL_LO 2711
`define SAVE_STATE_VGA_COL_HI 2720
`define SAVE_STATE_VGA_HS_CURR_STATE 2721
`define SAVE_STATE_VGA_VS_CURR_STATE 2722
`define SAVE_STATE_PPU_MEM_PAL_RAM_LO 2723
`define SAVE_STATE_PPU_MEM_PAL_RAM_HI 2754
`define SAVE_STATE_PPU_MEM_OAM_LO 2755
`define SAVE_STATE_PPU_MEM_OAM_HI 3010
`define SAVE_STATE_PPU_MEM_VRAM_LO 3011
`define SAVE_STATE_PPU_MEM_VRAM_HI 5058
`define SAVE_STATE_TRI_LEN_HALT 5059
`define SAVE_STATE_TRI_LIN_LOAD 5060
`define SAVE_STATE_TRI_LEN_LOAD 5061
`define SAVE_STATE_TRI_LIN_DATA 5062
`define SAVE_STATE_TRI_LEN_DATA 5063
`define SAVE_STATE_TRI_TIMER_PERIOD 5064
`define SAVE_STATE_TRI_SEQ_I 5065
`define SAVE_STATE_TRI_TIMER_COUNT 5066
`define SAVE_STATE_TRI_LIN_COUNT 5067
`define SAVE_STATE_TRI_LEN_COUNT 5068
`define SAVE_STATE_PUL_ENV_LOAD 5069
`define SAVE_STATE__SWEEP_LOAD 5070
`define SAVE_STATE__SWEEP_SIGS 5071
`define SAVE_STATE__DUTY 5072
`define SAVE_STATE__LEN_HALT 5073
`define SAVE_STATE__CONST_VOL 5074
`define SAVE_STATE__VOLUME 5075
`define SAVE_STATE__TIMER_PERIOD 5076
`define SAVE_STATE__LEN_LOAD 5077
`define SAVE_STATE__LEN_DATA 5078
`define SAVE_STATE__SEQ_I 5079
`define SAVE_STATE__TIMER_COUNT 5080
