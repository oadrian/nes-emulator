`default_nettype none
`include "ppu_defines.vh"


module sp_pixel (
    input clk, // Clock Enable (PPU Clock = Master clock/4)
    input rst_n  // Asynchronous reset active low
);

endmodule