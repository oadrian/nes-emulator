
`define SAVE_STATE_BITS ($clog2(4432))

`define SAVE_STATE_LAST_ADDRESS 4432

`define SAVE_STATE_CPU_UCODE_INDEX 0
`define SAVE_STATE_CPU_INSTR_CTRL_INDEX 1
`define SAVE_STATE_CPU_STATE 2
`define SAVE_STATE_CPU_NMI_ACTIVE 3
`define SAVE_STATE_CPU_RESET_ACTIVE 4
`define SAVE_STATE_CPU_CURRENT_INTERRUPT 5
`define SAVE_STATE_CPU_A 6
`define SAVE_STATE_CPU_X 7
`define SAVE_STATE_CPU_Y 8
`define SAVE_STATE_CPU_SP 9
`define SAVE_STATE_CPU_N_FLAG 10
`define SAVE_STATE_CPU_V_FLAG 11
`define SAVE_STATE_CPU_D_FLAG 12
`define SAVE_STATE_CPU_I_FLAG 13
`define SAVE_STATE_CPU_Z_FLAG 14
`define SAVE_STATE_CPU_C_FLAG 15
`define SAVE_STATE_CPU_PC 16
`define SAVE_STATE_CPU_R_DATA_BUFFER 17
`define SAVE_STATE_CPU_ADDR 18
`define SAVE_STATE_CPU_ALU_OUT 19
`define SAVE_STATE_CPU_ALU_C_OUT 20
`define SAVE_STATE_CPU_ALU_V_OUT 21
`define SAVE_STATE_CPU_ALU_Z_OUT 22
`define SAVE_STATE_CPU_ALU_N_OUT 23
`define SAVE_STATE_CPU_MEM_CPU_RAM_LO 24
`define SAVE_STATE_CPU_MEM_CPU_RAM_HI 2071
`define SAVE_STATE_CPU_MEM_READ_DATA 2072
`define SAVE_STATE_CPU_MEM_PREV_REG_EN 2073
`define SAVE_STATE_CPU_MEM_PREV_BUT_RD 2074
`define SAVE_STATE_CPU_MEM_PREV_APU_RD 2075
`define SAVE_STATE_PPU_PPUCTRL_OUT 2076
`define SAVE_STATE_PPU_PPUMASK_OUT 2077
`define SAVE_STATE_PPU_OAMDMA_OUT 2078
`define SAVE_STATE_PPU_OAMADDR_OUT 2079
`define SAVE_STATE_PPU_WR_CURR_STATE 2080
`define SAVE_STATE_PPU_REG_DATA_OUT 2081
`define SAVE_STATE_PPU_READ_BUF_CURR 2082
`define SAVE_STATE_PPU_PPUSTATUS_OUT 2083
`define SAVE_STATE_PPU_FORCE_VBLANK_CLR0 2084
`define SAVE_STATE_PPU_FORCE_VBLANK_CLR1 2085
`define SAVE_STATE_PPU_FX 2086
`define SAVE_STATE_PPU_TADDR  2087
`define SAVE_STATE_PPU_VADDR 2088
`define SAVE_STATE_VGA_ROW 2089
`define SAVE_STATE_VGA_COL 2090
`define SAVE_STATE_VGA_HS_CURR_STATE 2091
`define SAVE_STATE_VGA_VS_CURR_STATE 2092
`define SAVE_STATE_PPU_ROW 2093
`define SAVE_STATE_PPU_COL 2094
`define SAVE_STATE_PPU_HS_CURR_STATE 2095
`define SAVE_STATE_PPU_VS_CURR_STATE 2096
`define SAVE_STATE_PPU_MEM_PAL_RAM_LO 2097
`define SAVE_STATE_PPU_MEM_PAL_RAM_HI 2128
`define SAVE_STATE_PPU_MEM_OAM_LO 2129
`define SAVE_STATE_PPU_MEM_OAM_HI 2384
`define SAVE_STATE_PPU_MEM_VRAM_LO 2385
`define SAVE_STATE_PPU_MEM_VRAM_HI 4432
