`default_nettype none

module frame_counter (
  input logic clk, rst_l,
  input logic cpu_clock_en,
  
  output logic interrupt,
  output logic quarter_en, half_en);

  
endmodule: frame_counter
