
`define SAVE_STATE_BITS ($clog2(2072))

`define SAVE_STATE_LAST_ADDRESS 2072

`define SAVE_STATE_CPU_UCODE_INDEX 0
`define SAVE_STATE_CPU_INSTR_CTRL_INDEX 1
`define SAVE_STATE_CPU_STATE 2
`define SAVE_STATE_CPU_NMI_ACTIVE 3
`define SAVE_STATE_CPU_RESET_ACTIVE 4
`define SAVE_STATE_CPU_CURRENT_INTERUPT 5
`define SAVE_STATE_CPU_A 6
`define SAVE_STATE_CPU_X 7
`define SAVE_STATE_CPU_Y 8
`define SAVE_STATE_CPU_SP 9
`define SAVE_STATE_CPU_N_FLAG 10
`define SAVE_STATE_CPU_V_FLAG 11
`define SAVE_STATE_CPU_D_FLAG 12
`define SAVE_STATE_CPU_I_FLAG 13
`define SAVE_STATE_CPU_Z_FLAG 14
`define SAVE_STATE_CPU_C_FLAG 15
`define SAVE_STATE_CPU_PC 16
`define SAVE_STATE_CPU_R_DATA_BUFFER 17
`define SAVE_STATE_CPU_ADDR 18
`define SAVE_STATE_CPU_ALU_OUT 19
`define SAVE_STATE_CPU_ALU_C_OUT 20
`define SAVE_STATE_CPU_ALU_V_OUT 21
`define SAVE_STATE_CPU_ALU_Z_OUT 22
`define SAVE_STATE_CPU_ALU_N_OUT 23
`define SAVE_STATE_MEM_RAM_LO 24
`define SAVE_STATE_MEM_RAM_HI 2071
`define SAVE_STATE_MEM_READ_DATA 2072
