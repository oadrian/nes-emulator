`default_nettype none

module mixer(
    input  logic [3:0] pulse1, pulse2, triangle, noise,
    input  logic [6:0] dmc,
    output logic [15:0] out);

    logic [0:30][15:0] pulse_table;
    logic [0:202][15:0] tnd_table;
    logic [15:0] pulse_out, tnd_out, unsigned_out;

    assign pulse_out = pulse_table[pulse1 + pulse2];
    assign tnd_out = tnd_table[3*triangle + 2*noise + dmc];

    assign unsigned_out = pulse_out + tnd_out;
    assign out = {~unsigned_out[15], unsigned_out[14:0]};

    assign pulse_table = {
    16'd00000, 16'd00760, 16'd01503, 16'd02228, 16'd02936, 16'd03627, 16'd04303, 16'd04963, 
    16'd05609, 16'd06240, 16'd06857, 16'd07461, 16'd08053, 16'd08631, 16'd09198, 16'd09752, 
    16'd10295, 16'd10828, 16'd11349, 16'd11860, 16'd12361, 16'd12852, 16'd13334, 16'd13806, 
    16'd14270, 16'd14725, 16'd15171, 16'd15609, 16'd16039, 16'd16461, 16'd16876
    };

    assign tnd_table = {
    16'd00000, 16'd00439, 16'd00874, 16'd01306, 16'd01734, 16'd02159, 16'd02581, 16'd02999, 
    16'd03414, 16'd03826, 16'd04234, 16'd04639, 16'd05041, 16'd05440, 16'd05836, 16'd06229, 
    16'd06618, 16'd07005, 16'd07389, 16'd07769, 16'd08147, 16'd08522, 16'd08894, 16'd09264, 
    16'd09630, 16'd09994, 16'd10356, 16'd10714, 16'd11070, 16'd11423, 16'd11774, 16'd12122, 
    16'd12468, 16'd12811, 16'd13151, 16'd13490, 16'd13825, 16'd14159, 16'd14490, 16'd14818, 
    16'd15145, 16'd15469, 16'd15790, 16'd16110, 16'd16427, 16'd16742, 16'd17055, 16'd17366, 
    16'd17674, 16'd17981, 16'd18285, 16'd18588, 16'd18888, 16'd19186, 16'd19483, 16'd19777, 
    16'd20069, 16'd20359, 16'd20648, 16'd20934, 16'd21219, 16'd21502, 16'd21783, 16'd22062, 
    16'd22339, 16'd22614, 16'd22888, 16'd23160, 16'd23430, 16'd23699, 16'd23965, 16'd24230, 
    16'd24494, 16'd24755, 16'd25015, 16'd25274, 16'd25531, 16'd25786, 16'd26039, 16'd26291, 
    16'd26542, 16'd26791, 16'd27038, 16'd27284, 16'd27528, 16'd27771, 16'd28013, 16'd28253, 
    16'd28491, 16'd28728, 16'd28964, 16'd29198, 16'd29431, 16'd29662, 16'd29892, 16'd30121, 
    16'd30348, 16'd30574, 16'd30799, 16'd31022, 16'd31245, 16'd31465, 16'd31685, 16'd31903, 
    16'd32120, 16'd32336, 16'd32550, 16'd32764, 16'd32976, 16'd33187, 16'd33396, 16'd33605, 
    16'd33812, 16'd34018, 16'd34223, 16'd34427, 16'd34630, 16'd34831, 16'd35032, 16'd35231, 
    16'd35429, 16'd35627, 16'd35823, 16'd36018, 16'd36212, 16'd36405, 16'd36596, 16'd36787, 
    16'd36977, 16'd37166, 16'd37354, 16'd37540, 16'd37726, 16'd37911, 16'd38095, 16'd38278, 
    16'd38460, 16'd38640, 16'd38820, 16'd38999, 16'd39178, 16'd39355, 16'd39531, 16'd39706, 
    16'd39881, 16'd40054, 16'd40227, 16'd40399, 16'd40570, 16'd40740, 16'd40909, 16'd41077, 
    16'd41244, 16'd41411, 16'd41577, 16'd41742, 16'd41906, 16'd42069, 16'd42231, 16'd42393, 
    16'd42554, 16'd42714, 16'd42873, 16'd43032, 16'd43189, 16'd43346, 16'd43503, 16'd43658, 
    16'd43813, 16'd43966, 16'd44120, 16'd44272, 16'd44424, 16'd44575, 16'd44725, 16'd44874, 
    16'd45023, 16'd45171, 16'd45319, 16'd45465, 16'd45611, 16'd45757, 16'd45901, 16'd46045, 
    16'd46188, 16'd46331, 16'd46473, 16'd46614, 16'd46755, 16'd46895, 16'd47034, 16'd47173, 
    16'd47311, 16'd47448, 16'd47585, 16'd47721, 16'd47857, 16'd47992, 16'd48126, 16'd48260, 
    16'd48393, 16'd48525, 16'd48657
    };

endmodule : mixer